module StopWatchModule(/*AUTOARG*/);

   input i_clk;
   input i_rstn;
   input i_right;
   input i_left;
   input i_up;
   input i_down;

   
